`timescale 1ns/10ps
`define CYCLE   20.0   
`include "interface.sv"
`include "test.sv"
`include "LCD_CTRL.v"
